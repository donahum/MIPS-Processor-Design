/*
  Eric Villasenor
  evillase@gmail.com

  register file test bench
*/

// mapped needs this
`include "register_file_if.vh"

// mapped timing needs this. 1ns is too fast
`timescale 1 ns / 1 ns

module register_file_tb;

  parameter PERIOD = 10;

  logic CLK = 0, nRST;

  // test vars
  	//int v1 = 1;
  	//int v2 = 4721;
  	//int v3 = 25119;

  // clock
  always #(PERIOD/2) CLK++;

  // interface
  register_file_if rfif ();
  // test program
  test PROG (CLK, nRST, rfif);
  // DUT
`ifndef MAPPED
  register_file DUT(CLK, nRST, rfif);
`else
  register_file DUT(
    .\rfif.rdat2 (rfif.rdat2),
    .\rfif.rdat1 (rfif.rdat1),
    .\rfif.wdat (rfif.wdat),
    .\rfif.rsel2 (rfif.rsel2),
    .\rfif.rsel1 (rfif.rsel1),
    .\rfif.wsel (rfif.wsel),
    .\rfif.WEN (rfif.WEN),
    .\nRST (nRST),
    .\CLK (CLK)
  );
`endif

/*initial begin
	
end*/

task writeAndRead (input bit [4:0] wr_sel, [31:0] wr_dat);
	rfif.WEN = 0;
	rfif.wsel = '0;
	rfif.rsel1 = '0;
	rfif.rsel2 = '0;
	rfif.wdat = '0;
	#(PERIOD);

	rfif.WEN = 1;
	rfif.wsel = wr_sel;
	rfif.wdat = wr_dat;
	#(PERIOD);

	rfif.WEN = 0;
	rfif.wsel = '0;
	rfif.wdat = '0;
	rfif.rsel1 = wr_sel;
	rfif.rsel2 = wr_sel;
	#(PERIOD);

	rfif.WEN = 1;
	rfif.wsel = wr_sel;
	rfif.wdat = '0;
	#(PERIOD);

	rfif.WEN = 0;
	rfif.wsel = '0;
	rfif.rsel1 = '0;
	rfif.rsel2 = '0;
	rfif.wdat = '0;
	#(PERIOD);
endtask

endmodule

program test (
  input logic CLK,
  output logic nRST, register_file_if.tb tbrf
);
  parameter PERIOD = 10;
  initial begin
	$monitor("@%00g CLK = %b nRST = %b", $time, CLK, nRST);

	#(PERIOD);
	nRST = 1'b0;
	#(PERIOD);
	nRST = 1'b1;
    
	/*for(int i = 0; i < 32; i++)
	begin
		writeAndRead(i, 'hFFFFFFFF);
	end*/

	#(PERIOD);
	#(PERIOD);
	#(PERIOD);
	#(PERIOD);

	tbrf.WEN = 0;
	tbrf.wsel = '0;
	tbrf.rsel1 = '0;
	tbrf.rsel2 = '1;
	tbrf.wdat = '1;

	#(PERIOD);
	#(PERIOD);
	#(PERIOD);
	#(PERIOD);

	/*
	//test writing to reg1
	#(PERIOD);
	nRST = 1'b1;
	tbrf.WEN = 1'b1;
	tbrf.wsel = 5'b11111;
	tbrf.wdat = '1;
	#(PERIOD);

	//test writing to reg2
	#(PERIOD);
	nRST = 1'b1;
	tbrf.WEN = 1'b1;
	tbrf.wsel = 5'b11111;
	tbrf.wdat = '0;
	#(PERIOD);
	
	//check regs 1 and 2 to see if value held in one, not seen everywhere
	#(PERIOD);
	tbrf.WEN = 1'b0;
	tbrf.rsel1 = 5'b11111;
	tbrf.rsel2 = 5'b00010;
	#(PERIOD);
	
	//test async reset
	#(PERIOD);
	nRST = 1'b0;
	#(PERIOD);

	//test that values reset
	#(PERIOD);
	nRST = 1'b1;
	tbrf.rsel1 = 5'b00001;
	tbrf.rsel2 = 5'b11111;
	#(PERIOD);

	//test writing to reg0
	#(PERIOD);
	tbrf.WEN = 1'b1;
	tbrf.wsel = 5'b00000;
	tbrf.rsel1 = 5'b00000;
	tbrf.rsel2 = 5'b00001;
	#(PERIOD);*/

	//$finish;
  end
endprogram
